//-------------------------------------------------------------------------
//      test_memory.vhd                                                  --
//      Stephen Kempf                                                    --
//      Summer 2005                                                      --
//                                                                       --
//      Revised 3-15-2006                                                --
//              3-22-2007                                                --
//              7-26-2013                                                --
//                                                                       --
//      For use with ECE 385 Experment 6                                 --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------

// This memory has similar behavior to the SRAM IC on the DE2 board.  This
// file should be used for simulations only.  In simulation, this memory is
// guaranteed to work at least as well as the actual memory (that is, the
// actual memory may require more careful treatment than this test memory).

// To use, you should create a seperate top-level entity for simulation
// that connects this memory module to your computer.  You can create this
// extra entity either in the same project (temporarily setting it to be the
// top module) or in a new one, and create a new vector waveform file for it.


module test_memory ( input 			Clk,
							input          Reset, 
                     inout  [15:0]  I_O,
                     input  [19:0]  A,
                     input          CE,
                                    UB,
                                    LB,
                                    OE,
                                    WE );
												
   parameter size = 2000; // expand memory as needed (current is 64 words)
	 
   logic [15:0] mem_array [size-1:0];
   logic [15:0] mem_out;
   logic [15:0] I_O_wire;
	 
   assign mem_out = mem_array[A[19:0]];  //ATTENTION: Size here must correspond to size of
              // memory vector above.  Current size is 64, so the slice must be 6 bits.  If size were 1024,
              // slice would have to be 10 bits.  (There are three more places below where values must stay
              // consistent as well.)
	 
   always_comb
   begin
      I_O_wire = 16'bZZZZZZZZZZZZZZZZ;

      if (~CE && ~OE && WE) begin
         if (~UB)
            I_O_wire[15:8] = mem_out[15:8];
				
         if (~LB)
            I_O_wire[7:0] = mem_out[7:0];
		end
   end
	  
   always_ff @ (posedge Clk or posedge Reset)
   begin
		if(Reset)   // Insert initial memory contents here
		begin
mem_array[ 0 ] <= 16'h0;
mem_array[ 1 ] <= 16'h0;
mem_array[ 2 ] <= 16'h0;
mem_array[ 3 ] <= 16'h0;
mem_array[ 4 ] <= 16'h0;
mem_array[ 5 ] <= 16'h0;
mem_array[ 6 ] <= 16'h0;
mem_array[ 7 ] <= 16'h0;
mem_array[ 8 ] <= 16'h0;
mem_array[ 9 ] <= 16'h0;
mem_array[ 10 ] <= 16'h0;
mem_array[ 11 ] <= 16'h0;
mem_array[ 12 ] <= 16'h0;
mem_array[ 13 ] <= 16'h0;
mem_array[ 14 ] <= 16'h0;
mem_array[ 15 ] <= 16'h0;
mem_array[ 16 ] <= 16'h7bdf;
mem_array[ 17 ] <= 16'h0;
mem_array[ 18 ] <= 16'h0;
mem_array[ 19 ] <= 16'h0;
mem_array[ 20 ] <= 16'h0;
mem_array[ 21 ] <= 16'h0;
mem_array[ 22 ] <= 16'h0;
mem_array[ 23 ] <= 16'h0;
mem_array[ 24 ] <= 16'h0;
mem_array[ 25 ] <= 16'h0;
mem_array[ 26 ] <= 16'h0;
mem_array[ 27 ] <= 16'h0;
mem_array[ 28 ] <= 16'h0;
mem_array[ 29 ] <= 16'h0;
mem_array[ 30 ] <= 16'h0;
mem_array[ 31 ] <= 16'h0;
mem_array[ 32 ] <= 16'h0;
mem_array[ 33 ] <= 16'h0;
mem_array[ 34 ] <= 16'h0;
mem_array[ 35 ] <= 16'h0;
mem_array[ 36 ] <= 16'h0;
mem_array[ 37 ] <= 16'h0;
mem_array[ 38 ] <= 16'h0;
mem_array[ 39 ] <= 16'h0;
mem_array[ 40 ] <= 16'h0;
mem_array[ 41 ] <= 16'h0;
mem_array[ 42 ] <= 16'h1;
mem_array[ 43 ] <= 16'h1;
mem_array[ 44 ] <= 16'h1;
mem_array[ 45 ] <= 16'h1;
mem_array[ 46 ] <= 16'h1;
mem_array[ 47 ] <= 16'h1;
mem_array[ 48 ] <= 16'h1;
mem_array[ 49 ] <= 16'h1;
mem_array[ 50 ] <= 16'h1;
mem_array[ 51 ] <= 16'h1;
mem_array[ 52 ] <= 16'h1;
mem_array[ 53 ] <= 16'h1;
mem_array[ 54 ] <= 16'h0;
mem_array[ 55 ] <= 16'h0;
mem_array[ 56 ] <= 16'h0;
mem_array[ 57 ] <= 16'h0;
mem_array[ 58 ] <= 16'h0;
mem_array[ 59 ] <= 16'h0;
mem_array[ 60 ] <= 16'h0;
mem_array[ 61 ] <= 16'h0;
mem_array[ 62 ] <= 16'h0;
mem_array[ 63 ] <= 16'h0;
mem_array[ 64 ] <= 16'h0;
mem_array[ 65 ] <= 16'h0;
mem_array[ 66 ] <= 16'h0;
mem_array[ 67 ] <= 16'h0;
mem_array[ 68 ] <= 16'h0;
mem_array[ 69 ] <= 16'h0;
mem_array[ 70 ] <= 16'h0;
mem_array[ 71 ] <= 16'h0;
mem_array[ 72 ] <= 16'h1;
mem_array[ 73 ] <= 16'h1;
mem_array[ 74 ] <= 16'h1;
mem_array[ 75 ] <= 16'hb241;
mem_array[ 76 ] <= 16'hb241;
mem_array[ 77 ] <= 16'hb241;
mem_array[ 78 ] <= 16'hb241;
mem_array[ 79 ] <= 16'h1;
mem_array[ 80 ] <= 16'hb241;
mem_array[ 81 ] <= 16'h9981;
mem_array[ 82 ] <= 16'h9981;
mem_array[ 83 ] <= 16'h9981;
mem_array[ 84 ] <= 16'h9981;
mem_array[ 85 ] <= 16'h1;
mem_array[ 86 ] <= 16'h1;
mem_array[ 87 ] <= 16'h1;
mem_array[ 88 ] <= 16'h0;
mem_array[ 89 ] <= 16'h0;
mem_array[ 90 ] <= 16'h0;
mem_array[ 91 ] <= 16'h0;
mem_array[ 92 ] <= 16'h0;
mem_array[ 93 ] <= 16'h0;
mem_array[ 94 ] <= 16'h0;
mem_array[ 95 ] <= 16'h0;
mem_array[ 96 ] <= 16'h0;
mem_array[ 97 ] <= 16'h0;
mem_array[ 98 ] <= 16'h0;
mem_array[ 99 ] <= 16'h0;
mem_array[ 100 ] <= 16'h0;
mem_array[ 101 ] <= 16'h0;
mem_array[ 102 ] <= 16'h0;
mem_array[ 103 ] <= 16'h1;
mem_array[ 104 ] <= 16'h1;
mem_array[ 105 ] <= 16'hb241;
mem_array[ 106 ] <= 16'hb241;
mem_array[ 107 ] <= 16'hb241;
mem_array[ 108 ] <= 16'hb241;
mem_array[ 109 ] <= 16'hb241;
mem_array[ 110 ] <= 16'hb241;
mem_array[ 111 ] <= 16'h1;
mem_array[ 112 ] <= 16'hb241;
mem_array[ 113 ] <= 16'hb241;
mem_array[ 114 ] <= 16'hb241;
mem_array[ 115 ] <= 16'hb241;
mem_array[ 116 ] <= 16'h9981;
mem_array[ 117 ] <= 16'h9981;
mem_array[ 118 ] <= 16'h9981;
mem_array[ 119 ] <= 16'h1;
mem_array[ 120 ] <= 16'h1;
mem_array[ 121 ] <= 16'h0;
mem_array[ 122 ] <= 16'h0;
mem_array[ 123 ] <= 16'h0;
mem_array[ 124 ] <= 16'h0;
mem_array[ 125 ] <= 16'h0;
mem_array[ 126 ] <= 16'h0;
mem_array[ 127 ] <= 16'h0;
mem_array[ 128 ] <= 16'h0;
mem_array[ 129 ] <= 16'h0;
mem_array[ 130 ] <= 16'h0;
mem_array[ 131 ] <= 16'h0;
mem_array[ 132 ] <= 16'h0;
mem_array[ 133 ] <= 16'h1;
mem_array[ 134 ] <= 16'h1;
mem_array[ 135 ] <= 16'hcb01;
mem_array[ 136 ] <= 16'hcb01;
mem_array[ 137 ] <= 16'hcb01;
mem_array[ 138 ] <= 16'hcb01;
mem_array[ 139 ] <= 16'hcb01;
mem_array[ 140 ] <= 16'hcb01;
mem_array[ 141 ] <= 16'hcb01;
mem_array[ 142 ] <= 16'h1;
mem_array[ 143 ] <= 16'h1;
mem_array[ 144 ] <= 16'hb241;
mem_array[ 145 ] <= 16'hb241;
mem_array[ 146 ] <= 16'hb241;
mem_array[ 147 ] <= 16'hb241;
mem_array[ 148 ] <= 16'hb241;
mem_array[ 149 ] <= 16'hb241;
mem_array[ 150 ] <= 16'h9981;
mem_array[ 151 ] <= 16'h9981;
mem_array[ 152 ] <= 16'h9981;
mem_array[ 153 ] <= 16'h1;
mem_array[ 154 ] <= 16'h6b5b;
mem_array[ 155 ] <= 16'h0;
mem_array[ 156 ] <= 16'h0;
mem_array[ 157 ] <= 16'h0;
mem_array[ 158 ] <= 16'h0;
mem_array[ 159 ] <= 16'h0;
mem_array[ 160 ] <= 16'h0;
mem_array[ 161 ] <= 16'h0;
mem_array[ 162 ] <= 16'h0;
mem_array[ 163 ] <= 16'h0;
mem_array[ 164 ] <= 16'h1;
mem_array[ 165 ] <= 16'h1;
mem_array[ 166 ] <= 16'hcb01;
mem_array[ 167 ] <= 16'hcb01;
mem_array[ 168 ] <= 16'hcb01;
mem_array[ 169 ] <= 16'hcb01;
mem_array[ 170 ] <= 16'hcb01;
mem_array[ 171 ] <= 16'hb241;
mem_array[ 172 ] <= 16'hcb01;
mem_array[ 173 ] <= 16'hcb01;
mem_array[ 174 ] <= 16'h1;
mem_array[ 175 ] <= 16'h4901;
mem_array[ 176 ] <= 16'hcb01;
mem_array[ 177 ] <= 16'hb241;
mem_array[ 178 ] <= 16'hb241;
mem_array[ 179 ] <= 16'hb241;
mem_array[ 180 ] <= 16'hb241;
mem_array[ 181 ] <= 16'hb241;
mem_array[ 182 ] <= 16'hb241;
mem_array[ 183 ] <= 16'h9981;
mem_array[ 184 ] <= 16'h9981;
mem_array[ 185 ] <= 16'h9981;
mem_array[ 186 ] <= 16'h1;
mem_array[ 187 ] <= 16'h9ce7;
mem_array[ 188 ] <= 16'h0;
mem_array[ 189 ] <= 16'h0;
mem_array[ 190 ] <= 16'h0;
mem_array[ 191 ] <= 16'h0;
mem_array[ 192 ] <= 16'h0;
mem_array[ 193 ] <= 16'h0;
mem_array[ 194 ] <= 16'h0;
mem_array[ 195 ] <= 16'h0;
mem_array[ 196 ] <= 16'h1;
mem_array[ 197 ] <= 16'h1;
mem_array[ 198 ] <= 16'hcb01;
mem_array[ 199 ] <= 16'hb241;
mem_array[ 200 ] <= 16'hcb01;
mem_array[ 201 ] <= 16'hcb01;
mem_array[ 202 ] <= 16'hcb01;
mem_array[ 203 ] <= 16'hcb01;
mem_array[ 204 ] <= 16'hcb01;
mem_array[ 205 ] <= 16'hcb01;
mem_array[ 206 ] <= 16'h1;
mem_array[ 207 ] <= 16'hcb01;
mem_array[ 208 ] <= 16'hcb01;
mem_array[ 209 ] <= 16'hcb01;
mem_array[ 210 ] <= 16'hcb01;
mem_array[ 211 ] <= 16'hb241;
mem_array[ 212 ] <= 16'hb241;
mem_array[ 213 ] <= 16'hb241;
mem_array[ 214 ] <= 16'hb241;
mem_array[ 215 ] <= 16'hb241;
mem_array[ 216 ] <= 16'h9981;
mem_array[ 217 ] <= 16'h9981;
mem_array[ 218 ] <= 16'h9981;
mem_array[ 219 ] <= 16'h1;
mem_array[ 220 ] <= 16'h0;
mem_array[ 221 ] <= 16'h0;
mem_array[ 222 ] <= 16'h0;
mem_array[ 223 ] <= 16'h0;
mem_array[ 224 ] <= 16'h0;
mem_array[ 225 ] <= 16'h0;
mem_array[ 226 ] <= 16'h0;
mem_array[ 227 ] <= 16'h1;
mem_array[ 228 ] <= 16'hcb01;
mem_array[ 229 ] <= 16'h1;
mem_array[ 230 ] <= 16'hcb01;
mem_array[ 231 ] <= 16'hb241;
mem_array[ 232 ] <= 16'hcb01;
mem_array[ 233 ] <= 16'hba81;
mem_array[ 234 ] <= 16'hcb01;
mem_array[ 235 ] <= 16'hcb01;
mem_array[ 236 ] <= 16'hcb01;
mem_array[ 237 ] <= 16'hcb01;
mem_array[ 238 ] <= 16'h1;
mem_array[ 239 ] <= 16'hcb01;
mem_array[ 240 ] <= 16'hcb01;
mem_array[ 241 ] <= 16'hcb01;
mem_array[ 242 ] <= 16'hcb01;
mem_array[ 243 ] <= 16'hcb01;
mem_array[ 244 ] <= 16'hb241;
mem_array[ 245 ] <= 16'hb241;
mem_array[ 246 ] <= 16'hb241;
mem_array[ 247 ] <= 16'hb241;
mem_array[ 248 ] <= 16'hb241;
mem_array[ 249 ] <= 16'h9981;
mem_array[ 250 ] <= 16'h9981;
mem_array[ 251 ] <= 16'h1;
mem_array[ 252 ] <= 16'h1;
mem_array[ 253 ] <= 16'h0;
mem_array[ 254 ] <= 16'h0;
mem_array[ 255 ] <= 16'h0;
mem_array[ 256 ] <= 16'h0;
mem_array[ 257 ] <= 16'h0;
mem_array[ 258 ] <= 16'h1;
mem_array[ 259 ] <= 16'h1;
mem_array[ 260 ] <= 16'hcb01;
mem_array[ 261 ] <= 16'h1;
mem_array[ 262 ] <= 16'hcb01;
mem_array[ 263 ] <= 16'hcb01;
mem_array[ 264 ] <= 16'hcb01;
mem_array[ 265 ] <= 16'hcb01;
mem_array[ 266 ] <= 16'hcb01;
mem_array[ 267 ] <= 16'hcb01;
mem_array[ 268 ] <= 16'hb241;
mem_array[ 269 ] <= 16'h1;
mem_array[ 270 ] <= 16'h1;
mem_array[ 271 ] <= 16'hcb01;
mem_array[ 272 ] <= 16'hcb01;
mem_array[ 273 ] <= 16'hcb01;
mem_array[ 274 ] <= 16'hcb01;
mem_array[ 275 ] <= 16'hcb01;
mem_array[ 276 ] <= 16'hcb01;
mem_array[ 277 ] <= 16'hb241;
mem_array[ 278 ] <= 16'hb241;
mem_array[ 279 ] <= 16'hb241;
mem_array[ 280 ] <= 16'hb241;
mem_array[ 281 ] <= 16'hb241;
mem_array[ 282 ] <= 16'h9981;
mem_array[ 283 ] <= 16'h1;
mem_array[ 284 ] <= 16'h1;
mem_array[ 285 ] <= 16'h1;
mem_array[ 286 ] <= 16'h0;
mem_array[ 287 ] <= 16'h0;
mem_array[ 288 ] <= 16'h0;
mem_array[ 289 ] <= 16'h0;
mem_array[ 290 ] <= 16'h1;
mem_array[ 291 ] <= 16'hcb01;
mem_array[ 292 ] <= 16'hdbc5;
mem_array[ 293 ] <= 16'h1;
mem_array[ 294 ] <= 16'hdbc5;
mem_array[ 295 ] <= 16'hdbc5;
mem_array[ 296 ] <= 16'hdbc5;
mem_array[ 297 ] <= 16'hdbc5;
mem_array[ 298 ] <= 16'hcb41;
mem_array[ 299 ] <= 16'hcb01;
mem_array[ 300 ] <= 16'hcb01;
mem_array[ 301 ] <= 16'h1;
mem_array[ 302 ] <= 16'hcb01;
mem_array[ 303 ] <= 16'hcb01;
mem_array[ 304 ] <= 16'hcb01;
mem_array[ 305 ] <= 16'hcb01;
mem_array[ 306 ] <= 16'hcb01;
mem_array[ 307 ] <= 16'hcb01;
mem_array[ 308 ] <= 16'hcb01;
mem_array[ 309 ] <= 16'hcb01;
mem_array[ 310 ] <= 16'hb241;
mem_array[ 311 ] <= 16'hb241;
mem_array[ 312 ] <= 16'hb241;
mem_array[ 313 ] <= 16'hb241;
mem_array[ 314 ] <= 16'hb241;
mem_array[ 315 ] <= 16'h1;
mem_array[ 316 ] <= 16'h9981;
mem_array[ 317 ] <= 16'h1;
mem_array[ 318 ] <= 16'h0;
mem_array[ 319 ] <= 16'h0;
mem_array[ 320 ] <= 16'h0;
mem_array[ 321 ] <= 16'h1;
mem_array[ 322 ] <= 16'h1;
mem_array[ 323 ] <= 16'hdbc5;
mem_array[ 324 ] <= 16'hdbc5;
mem_array[ 325 ] <= 16'h1;
mem_array[ 326 ] <= 16'h1;
mem_array[ 327 ] <= 16'hdbc5;
mem_array[ 328 ] <= 16'hdbc5;
mem_array[ 329 ] <= 16'hdbc5;
mem_array[ 330 ] <= 16'hdbc5;
mem_array[ 331 ] <= 16'hdbc5;
mem_array[ 332 ] <= 16'hcb01;
mem_array[ 333 ] <= 16'h1;
mem_array[ 334 ] <= 16'hcb01;
mem_array[ 335 ] <= 16'hcb01;
mem_array[ 336 ] <= 16'hcb01;
mem_array[ 337 ] <= 16'hcb01;
mem_array[ 338 ] <= 16'hcb01;
mem_array[ 339 ] <= 16'hcb01;
mem_array[ 340 ] <= 16'hcb01;
mem_array[ 341 ] <= 16'hcb01;
mem_array[ 342 ] <= 16'hb241;
mem_array[ 343 ] <= 16'hb241;
mem_array[ 344 ] <= 16'hb241;
mem_array[ 345 ] <= 16'hb241;
mem_array[ 346 ] <= 16'h1;
mem_array[ 347 ] <= 16'h9981;
mem_array[ 348 ] <= 16'h9981;
mem_array[ 349 ] <= 16'h1;
mem_array[ 350 ] <= 16'h1;
mem_array[ 351 ] <= 16'h0;
mem_array[ 352 ] <= 16'h0;
mem_array[ 353 ] <= 16'h1;
mem_array[ 354 ] <= 16'hdbc5;
mem_array[ 355 ] <= 16'hdbc5;
mem_array[ 356 ] <= 16'hdbc5;
mem_array[ 357 ] <= 16'hdbc5;
mem_array[ 358 ] <= 16'h1;
mem_array[ 359 ] <= 16'hdbc5;
mem_array[ 360 ] <= 16'hdbc5;
mem_array[ 361 ] <= 16'hcb01;
mem_array[ 362 ] <= 16'hdbc5;
mem_array[ 363 ] <= 16'hdbc5;
mem_array[ 364 ] <= 16'h7a03;
mem_array[ 365 ] <= 16'h1;
mem_array[ 366 ] <= 16'hcb01;
mem_array[ 367 ] <= 16'hcb01;
mem_array[ 368 ] <= 16'hcb01;
mem_array[ 369 ] <= 16'hcb01;
mem_array[ 370 ] <= 16'hcb01;
mem_array[ 371 ] <= 16'hcb01;
mem_array[ 372 ] <= 16'hcb01;
mem_array[ 373 ] <= 16'hcb01;
mem_array[ 374 ] <= 16'hcb01;
mem_array[ 375 ] <= 16'hb241;
mem_array[ 376 ] <= 16'hb241;
mem_array[ 377 ] <= 16'h1;
mem_array[ 378 ] <= 16'h1;
mem_array[ 379 ] <= 16'hb241;
mem_array[ 380 ] <= 16'h9981;
mem_array[ 381 ] <= 16'h9981;
mem_array[ 382 ] <= 16'h1;
mem_array[ 383 ] <= 16'h0;
mem_array[ 384 ] <= 16'h0;
mem_array[ 385 ] <= 16'h1;
mem_array[ 386 ] <= 16'hdbc5;
mem_array[ 387 ] <= 16'hdbc5;
mem_array[ 388 ] <= 16'hec07;
mem_array[ 389 ] <= 16'hf449;
mem_array[ 390 ] <= 16'h1;
mem_array[ 391 ] <= 16'h1;
mem_array[ 392 ] <= 16'hdbc5;
mem_array[ 393 ] <= 16'hdbc5;
mem_array[ 394 ] <= 16'hcb01;
mem_array[ 395 ] <= 16'hdbc5;
mem_array[ 396 ] <= 16'h1;
mem_array[ 397 ] <= 16'hcb01;
mem_array[ 398 ] <= 16'hcb01;
mem_array[ 399 ] <= 16'hcb01;
mem_array[ 400 ] <= 16'hcb01;
mem_array[ 401 ] <= 16'hcb01;
mem_array[ 402 ] <= 16'hcb01;
mem_array[ 403 ] <= 16'hcb01;
mem_array[ 404 ] <= 16'hcb01;
mem_array[ 405 ] <= 16'hcb01;
mem_array[ 406 ] <= 16'hcb01;
mem_array[ 407 ] <= 16'hb241;
mem_array[ 408 ] <= 16'h1;
mem_array[ 409 ] <= 16'h1;
mem_array[ 410 ] <= 16'hb241;
mem_array[ 411 ] <= 16'hb241;
mem_array[ 412 ] <= 16'h9981;
mem_array[ 413 ] <= 16'h9981;
mem_array[ 414 ] <= 16'h1;
mem_array[ 415 ] <= 16'h0;
mem_array[ 416 ] <= 16'h1;
mem_array[ 417 ] <= 16'h1;
mem_array[ 418 ] <= 16'hdbc5;
mem_array[ 419 ] <= 16'hf449;
mem_array[ 420 ] <= 16'hf449;
mem_array[ 421 ] <= 16'hf449;
mem_array[ 422 ] <= 16'hf449;
mem_array[ 423 ] <= 16'h1;
mem_array[ 424 ] <= 16'h1;
mem_array[ 425 ] <= 16'hdbc5;
mem_array[ 426 ] <= 16'hcb01;
mem_array[ 427 ] <= 16'hdbc5;
mem_array[ 428 ] <= 16'h1;
mem_array[ 429 ] <= 16'hdbc5;
mem_array[ 430 ] <= 16'hcb01;
mem_array[ 431 ] <= 16'hcb01;
mem_array[ 432 ] <= 16'hcb01;
mem_array[ 433 ] <= 16'hcb01;
mem_array[ 434 ] <= 16'hcb01;
mem_array[ 435 ] <= 16'hcb01;
mem_array[ 436 ] <= 16'hcb01;
mem_array[ 437 ] <= 16'hcb01;
mem_array[ 438 ] <= 16'hcb01;
mem_array[ 439 ] <= 16'h1;
mem_array[ 440 ] <= 16'h1;
mem_array[ 441 ] <= 16'hb241;
mem_array[ 442 ] <= 16'hb241;
mem_array[ 443 ] <= 16'hb241;
mem_array[ 444 ] <= 16'h9981;
mem_array[ 445 ] <= 16'h9981;
mem_array[ 446 ] <= 16'h1;
mem_array[ 447 ] <= 16'h1;
mem_array[ 448 ] <= 16'h1;
mem_array[ 449 ] <= 16'h1;
mem_array[ 450 ] <= 16'hdbc5;
mem_array[ 451 ] <= 16'hf449;
mem_array[ 452 ] <= 16'hdbc5;
mem_array[ 453 ] <= 16'hf449;
mem_array[ 454 ] <= 16'hf449;
mem_array[ 455 ] <= 16'hf449;
mem_array[ 456 ] <= 16'h1;
mem_array[ 457 ] <= 16'h1;
mem_array[ 458 ] <= 16'hdbc5;
mem_array[ 459 ] <= 16'hdbc5;
mem_array[ 460 ] <= 16'h1;
mem_array[ 461 ] <= 16'hdbc5;
mem_array[ 462 ] <= 16'hcb01;
mem_array[ 463 ] <= 16'hcb01;
mem_array[ 464 ] <= 16'hcb01;
mem_array[ 465 ] <= 16'hcb01;
mem_array[ 466 ] <= 16'hcb01;
mem_array[ 467 ] <= 16'hcb01;
mem_array[ 468 ] <= 16'hcb01;
mem_array[ 469 ] <= 16'hcb01;
mem_array[ 470 ] <= 16'h1;
mem_array[ 471 ] <= 16'h1;
mem_array[ 472 ] <= 16'hb241;
mem_array[ 473 ] <= 16'hb241;
mem_array[ 474 ] <= 16'hb241;
mem_array[ 475 ] <= 16'hb241;
mem_array[ 476 ] <= 16'h9981;
mem_array[ 477 ] <= 16'h9981;
mem_array[ 478 ] <= 16'h1;
mem_array[ 479 ] <= 16'h1;
mem_array[ 480 ] <= 16'h1;
mem_array[ 481 ] <= 16'h1;
mem_array[ 482 ] <= 16'hf449;
mem_array[ 483 ] <= 16'hf449;
mem_array[ 484 ] <= 16'hf449;
mem_array[ 485 ] <= 16'hdbc5;
mem_array[ 486 ] <= 16'hdbc5;
mem_array[ 487 ] <= 16'hf449;
mem_array[ 488 ] <= 16'hf449;
mem_array[ 489 ] <= 16'h1;
mem_array[ 490 ] <= 16'h1;
mem_array[ 491 ] <= 16'h1;
mem_array[ 492 ] <= 16'h1;
mem_array[ 493 ] <= 16'hdbc5;
mem_array[ 494 ] <= 16'hcb01;
mem_array[ 495 ] <= 16'hcb01;
mem_array[ 496 ] <= 16'hcb01;
mem_array[ 497 ] <= 16'hcb01;
mem_array[ 498 ] <= 16'hcb01;
mem_array[ 499 ] <= 16'h1;
mem_array[ 500 ] <= 16'h1;
mem_array[ 501 ] <= 16'h1;
mem_array[ 502 ] <= 16'hcb01;
mem_array[ 503 ] <= 16'hcb01;
mem_array[ 504 ] <= 16'hb241;
mem_array[ 505 ] <= 16'hb241;
mem_array[ 506 ] <= 16'hb241;
mem_array[ 507 ] <= 16'hb241;
mem_array[ 508 ] <= 16'h9981;
mem_array[ 509 ] <= 16'h9981;
mem_array[ 510 ] <= 16'h1;
mem_array[ 511 ] <= 16'h1;
mem_array[ 512 ] <= 16'h1;
mem_array[ 513 ] <= 16'h1;
mem_array[ 514 ] <= 16'hf449;
mem_array[ 515 ] <= 16'hf449;
mem_array[ 516 ] <= 16'hdbc5;
mem_array[ 517 ] <= 16'hf449;
mem_array[ 518 ] <= 16'hf449;
mem_array[ 519 ] <= 16'hf449;
mem_array[ 520 ] <= 16'hdbc5;
mem_array[ 521 ] <= 16'hf449;
mem_array[ 522 ] <= 16'hdbc5;
mem_array[ 523 ] <= 16'h1;
mem_array[ 524 ] <= 16'h1;
mem_array[ 525 ] <= 16'h1;
mem_array[ 526 ] <= 16'h1;
mem_array[ 527 ] <= 16'h1;
mem_array[ 528 ] <= 16'h1;
mem_array[ 529 ] <= 16'h1;
mem_array[ 530 ] <= 16'h1;
mem_array[ 531 ] <= 16'h1;
mem_array[ 532 ] <= 16'hcb01;
mem_array[ 533 ] <= 16'hcb01;
mem_array[ 534 ] <= 16'hcb01;
mem_array[ 535 ] <= 16'hcb01;
mem_array[ 536 ] <= 16'hcb01;
mem_array[ 537 ] <= 16'hb241;
mem_array[ 538 ] <= 16'hb241;
mem_array[ 539 ] <= 16'hb241;
mem_array[ 540 ] <= 16'h9981;
mem_array[ 541 ] <= 16'h9981;
mem_array[ 542 ] <= 16'h1;
mem_array[ 543 ] <= 16'h1;
mem_array[ 544 ] <= 16'h1;
mem_array[ 545 ] <= 16'h1;
mem_array[ 546 ] <= 16'h1;
mem_array[ 547 ] <= 16'hf449;
mem_array[ 548 ] <= 16'hf449;
mem_array[ 549 ] <= 16'hf449;
mem_array[ 550 ] <= 16'hf449;
mem_array[ 551 ] <= 16'hf449;
mem_array[ 552 ] <= 16'hec49;
mem_array[ 553 ] <= 16'hf449;
mem_array[ 554 ] <= 16'hf449;
mem_array[ 555 ] <= 16'h1;
mem_array[ 556 ] <= 16'hdbc5;
mem_array[ 557 ] <= 16'hdbc5;
mem_array[ 558 ] <= 16'hdbc5;
mem_array[ 559 ] <= 16'hcb01;
mem_array[ 560 ] <= 16'hcb01;
mem_array[ 561 ] <= 16'hcb01;
mem_array[ 562 ] <= 16'hcb01;
mem_array[ 563 ] <= 16'hcb01;
mem_array[ 564 ] <= 16'hcb01;
mem_array[ 565 ] <= 16'hcb01;
mem_array[ 566 ] <= 16'hcb01;
mem_array[ 567 ] <= 16'hcb01;
mem_array[ 568 ] <= 16'hcb01;
mem_array[ 569 ] <= 16'hb241;
mem_array[ 570 ] <= 16'hb241;
mem_array[ 571 ] <= 16'hb241;
mem_array[ 572 ] <= 16'h9981;
mem_array[ 573 ] <= 16'h9981;
mem_array[ 574 ] <= 16'h1;
mem_array[ 575 ] <= 16'h1;
mem_array[ 576 ] <= 16'h39cf;
mem_array[ 577 ] <= 16'h1;
mem_array[ 578 ] <= 16'hdbc5;
mem_array[ 579 ] <= 16'h1;
mem_array[ 580 ] <= 16'hf449;
mem_array[ 581 ] <= 16'hf449;
mem_array[ 582 ] <= 16'hdbc5;
mem_array[ 583 ] <= 16'hf449;
mem_array[ 584 ] <= 16'hf449;
mem_array[ 585 ] <= 16'hf449;
mem_array[ 586 ] <= 16'hf449;
mem_array[ 587 ] <= 16'h1;
mem_array[ 588 ] <= 16'hdbc5;
mem_array[ 589 ] <= 16'hdbc5;
mem_array[ 590 ] <= 16'hdbc5;
mem_array[ 591 ] <= 16'hcb01;
mem_array[ 592 ] <= 16'hcb01;
mem_array[ 593 ] <= 16'hcb01;
mem_array[ 594 ] <= 16'hcb01;
mem_array[ 595 ] <= 16'hcb01;
mem_array[ 596 ] <= 16'hcb01;
mem_array[ 597 ] <= 16'hcb01;
mem_array[ 598 ] <= 16'hcb01;
mem_array[ 599 ] <= 16'hcb01;
mem_array[ 600 ] <= 16'hcb01;
mem_array[ 601 ] <= 16'hb241;
mem_array[ 602 ] <= 16'hb241;
mem_array[ 603 ] <= 16'hb241;
mem_array[ 604 ] <= 16'h9981;
mem_array[ 605 ] <= 16'h1;
mem_array[ 606 ] <= 16'h1;
mem_array[ 607 ] <= 16'h1;
mem_array[ 608 ] <= 16'h0;
mem_array[ 609 ] <= 16'h1;
mem_array[ 610 ] <= 16'hdbc5;
mem_array[ 611 ] <= 16'hf449;
mem_array[ 612 ] <= 16'h1;
mem_array[ 613 ] <= 16'h1;
mem_array[ 614 ] <= 16'hf449;
mem_array[ 615 ] <= 16'hf449;
mem_array[ 616 ] <= 16'hf449;
mem_array[ 617 ] <= 16'hf449;
mem_array[ 618 ] <= 16'h1;
mem_array[ 619 ] <= 16'h1;
mem_array[ 620 ] <= 16'hcb01;
mem_array[ 621 ] <= 16'hdbc5;
mem_array[ 622 ] <= 16'hdbc5;
mem_array[ 623 ] <= 16'hcb01;
mem_array[ 624 ] <= 16'hcb01;
mem_array[ 625 ] <= 16'hcb01;
mem_array[ 626 ] <= 16'hcb01;
mem_array[ 627 ] <= 16'hcb01;
mem_array[ 628 ] <= 16'hcb01;
mem_array[ 629 ] <= 16'hcb01;
mem_array[ 630 ] <= 16'hcb01;
mem_array[ 631 ] <= 16'hcb01;
mem_array[ 632 ] <= 16'hcb01;
mem_array[ 633 ] <= 16'hb241;
mem_array[ 634 ] <= 16'hb241;
mem_array[ 635 ] <= 16'hb241;
mem_array[ 636 ] <= 16'h9981;
mem_array[ 637 ] <= 16'h1;
mem_array[ 638 ] <= 16'h1;
mem_array[ 639 ] <= 16'h0;
mem_array[ 640 ] <= 16'h0;
mem_array[ 641 ] <= 16'h1;
mem_array[ 642 ] <= 16'hdbc5;
mem_array[ 643 ] <= 16'hdbc5;
mem_array[ 644 ] <= 16'hf449;
mem_array[ 645 ] <= 16'h1;
mem_array[ 646 ] <= 16'h1;
mem_array[ 647 ] <= 16'hf449;
mem_array[ 648 ] <= 16'hf449;
mem_array[ 649 ] <= 16'hf449;
mem_array[ 650 ] <= 16'h1;
mem_array[ 651 ] <= 16'h1;
mem_array[ 652 ] <= 16'hdbc5;
mem_array[ 653 ] <= 16'hdbc5;
mem_array[ 654 ] <= 16'hdbc5;
mem_array[ 655 ] <= 16'hcb01;
mem_array[ 656 ] <= 16'hcb01;
mem_array[ 657 ] <= 16'hcb01;
mem_array[ 658 ] <= 16'hcb01;
mem_array[ 659 ] <= 16'hcb01;
mem_array[ 660 ] <= 16'hcb01;
mem_array[ 661 ] <= 16'hcb01;
mem_array[ 662 ] <= 16'hcb01;
mem_array[ 663 ] <= 16'hcb01;
mem_array[ 664 ] <= 16'hcb01;
mem_array[ 665 ] <= 16'hb241;
mem_array[ 666 ] <= 16'hb241;
mem_array[ 667 ] <= 16'h801;
mem_array[ 668 ] <= 16'h1;
mem_array[ 669 ] <= 16'h9981;
mem_array[ 670 ] <= 16'h1;
mem_array[ 671 ] <= 16'h0;
mem_array[ 672 ] <= 16'h0;
mem_array[ 673 ] <= 16'h1;
mem_array[ 674 ] <= 16'h1;
mem_array[ 675 ] <= 16'hdbc5;
mem_array[ 676 ] <= 16'hf449;
mem_array[ 677 ] <= 16'hdbc5;
mem_array[ 678 ] <= 16'hf449;
mem_array[ 679 ] <= 16'h1;
mem_array[ 680 ] <= 16'h1;
mem_array[ 681 ] <= 16'h1;
mem_array[ 682 ] <= 16'h1;
mem_array[ 683 ] <= 16'hcb01;
mem_array[ 684 ] <= 16'hdbc5;
mem_array[ 685 ] <= 16'hcb01;
mem_array[ 686 ] <= 16'hdbc5;
mem_array[ 687 ] <= 16'hcb01;
mem_array[ 688 ] <= 16'hcb01;
mem_array[ 689 ] <= 16'hcb01;
mem_array[ 690 ] <= 16'hcb01;
mem_array[ 691 ] <= 16'hcb01;
mem_array[ 692 ] <= 16'hcb01;
mem_array[ 693 ] <= 16'hcb01;
mem_array[ 694 ] <= 16'hcb01;
mem_array[ 695 ] <= 16'hcb01;
mem_array[ 696 ] <= 16'hcb01;
mem_array[ 697 ] <= 16'hb241;
mem_array[ 698 ] <= 16'h1;
mem_array[ 699 ] <= 16'h1;
mem_array[ 700 ] <= 16'h9981;
mem_array[ 701 ] <= 16'h1001;
mem_array[ 702 ] <= 16'h1;
mem_array[ 703 ] <= 16'h0;
mem_array[ 704 ] <= 16'h0;
mem_array[ 705 ] <= 16'h0;
mem_array[ 706 ] <= 16'h1;
mem_array[ 707 ] <= 16'hdbc5;
mem_array[ 708 ] <= 16'hdbc5;
mem_array[ 709 ] <= 16'hf449;
mem_array[ 710 ] <= 16'hf449;
mem_array[ 711 ] <= 16'hf449;
mem_array[ 712 ] <= 16'hf449;
mem_array[ 713 ] <= 16'h1;
mem_array[ 714 ] <= 16'h1;
mem_array[ 715 ] <= 16'h1;
mem_array[ 716 ] <= 16'h1;
mem_array[ 717 ] <= 16'hdbc5;
mem_array[ 718 ] <= 16'hdbc5;
mem_array[ 719 ] <= 16'hcb01;
mem_array[ 720 ] <= 16'hcb01;
mem_array[ 721 ] <= 16'hcb01;
mem_array[ 722 ] <= 16'hcb01;
mem_array[ 723 ] <= 16'hcb01;
mem_array[ 724 ] <= 16'hcb01;
mem_array[ 725 ] <= 16'hcb01;
mem_array[ 726 ] <= 16'hcb01;
mem_array[ 727 ] <= 16'h71c1;
mem_array[ 728 ] <= 16'h1;
mem_array[ 729 ] <= 16'h1;
mem_array[ 730 ] <= 16'h1;
mem_array[ 731 ] <= 16'h9981;
mem_array[ 732 ] <= 16'h9981;
mem_array[ 733 ] <= 16'h1;
mem_array[ 734 ] <= 16'h0;
mem_array[ 735 ] <= 16'h0;
mem_array[ 736 ] <= 16'h0;
mem_array[ 737 ] <= 16'h0;
mem_array[ 738 ] <= 16'h1;
mem_array[ 739 ] <= 16'h1;
mem_array[ 740 ] <= 16'hdbc5;
mem_array[ 741 ] <= 16'hf449;
mem_array[ 742 ] <= 16'hdbc5;
mem_array[ 743 ] <= 16'hec49;
mem_array[ 744 ] <= 16'hf449;
mem_array[ 745 ] <= 16'hf449;
mem_array[ 746 ] <= 16'h1;
mem_array[ 747 ] <= 16'hdbc5;
mem_array[ 748 ] <= 16'h1;
mem_array[ 749 ] <= 16'h1;
mem_array[ 750 ] <= 16'h1;
mem_array[ 751 ] <= 16'h1;
mem_array[ 752 ] <= 16'h1;
mem_array[ 753 ] <= 16'h1;
mem_array[ 754 ] <= 16'h1;
mem_array[ 755 ] <= 16'h1;
mem_array[ 756 ] <= 16'h1;
mem_array[ 757 ] <= 16'h1;
mem_array[ 758 ] <= 16'h1;
mem_array[ 759 ] <= 16'h1;
mem_array[ 760 ] <= 16'hb241;
mem_array[ 761 ] <= 16'hb241;
mem_array[ 762 ] <= 16'hb241;
mem_array[ 763 ] <= 16'h9981;
mem_array[ 764 ] <= 16'h1;
mem_array[ 765 ] <= 16'h1;
mem_array[ 766 ] <= 16'h0;
mem_array[ 767 ] <= 16'h0;
mem_array[ 768 ] <= 16'h0;
mem_array[ 769 ] <= 16'h0;
mem_array[ 770 ] <= 16'h0;
mem_array[ 771 ] <= 16'h1;
mem_array[ 772 ] <= 16'hd383;
mem_array[ 773 ] <= 16'hdbc5;
mem_array[ 774 ] <= 16'hf449;
mem_array[ 775 ] <= 16'hf449;
mem_array[ 776 ] <= 16'hf449;
mem_array[ 777 ] <= 16'hf449;
mem_array[ 778 ] <= 16'h1;
mem_array[ 779 ] <= 16'hdbc5;
mem_array[ 780 ] <= 16'hdbc5;
mem_array[ 781 ] <= 16'hdbc5;
mem_array[ 782 ] <= 16'hcb01;
mem_array[ 783 ] <= 16'hcb01;
mem_array[ 784 ] <= 16'hcb01;
mem_array[ 785 ] <= 16'h30c1;
mem_array[ 786 ] <= 16'h1;
mem_array[ 787 ] <= 16'hcb01;
mem_array[ 788 ] <= 16'hcb01;
mem_array[ 789 ] <= 16'hcb01;
mem_array[ 790 ] <= 16'hcb01;
mem_array[ 791 ] <= 16'hcb01;
mem_array[ 792 ] <= 16'hb241;
mem_array[ 793 ] <= 16'hb241;
mem_array[ 794 ] <= 16'h99c1;
mem_array[ 795 ] <= 16'h9981;
mem_array[ 796 ] <= 16'h1;
mem_array[ 797 ] <= 16'h0;
mem_array[ 798 ] <= 16'h0;
mem_array[ 799 ] <= 16'h0;
mem_array[ 800 ] <= 16'h0;
mem_array[ 801 ] <= 16'h0;
mem_array[ 802 ] <= 16'h0;
mem_array[ 803 ] <= 16'h1;
mem_array[ 804 ] <= 16'h1;
mem_array[ 805 ] <= 16'hdbc5;
mem_array[ 806 ] <= 16'hcb01;
mem_array[ 807 ] <= 16'hdbc5;
mem_array[ 808 ] <= 16'hdbc5;
mem_array[ 809 ] <= 16'hdbc5;
mem_array[ 810 ] <= 16'h1;
mem_array[ 811 ] <= 16'hdbc5;
mem_array[ 812 ] <= 16'hdbc5;
mem_array[ 813 ] <= 16'hdbc5;
mem_array[ 814 ] <= 16'hcb01;
mem_array[ 815 ] <= 16'hcb01;
mem_array[ 816 ] <= 16'hcb01;
mem_array[ 817 ] <= 16'hcb01;
mem_array[ 818 ] <= 16'hcb01;
mem_array[ 819 ] <= 16'hcb01;
mem_array[ 820 ] <= 16'hcb01;
mem_array[ 821 ] <= 16'hcb01;
mem_array[ 822 ] <= 16'hcb01;
mem_array[ 823 ] <= 16'hb241;
mem_array[ 824 ] <= 16'hb241;
mem_array[ 825 ] <= 16'hb241;
mem_array[ 826 ] <= 16'h9981;
mem_array[ 827 ] <= 16'h1;
mem_array[ 828 ] <= 16'h0;
mem_array[ 829 ] <= 16'h0;
mem_array[ 830 ] <= 16'h0;
mem_array[ 831 ] <= 16'h0;
mem_array[ 832 ] <= 16'h0;
mem_array[ 833 ] <= 16'h0;
mem_array[ 834 ] <= 16'h0;
mem_array[ 835 ] <= 16'h0;
mem_array[ 836 ] <= 16'h1;
mem_array[ 837 ] <= 16'h1;
mem_array[ 838 ] <= 16'hdbc5;
mem_array[ 839 ] <= 16'h1;
mem_array[ 840 ] <= 16'h1;
mem_array[ 841 ] <= 16'h1;
mem_array[ 842 ] <= 16'h1;
mem_array[ 843 ] <= 16'h1;
mem_array[ 844 ] <= 16'h1;
mem_array[ 845 ] <= 16'h1;
mem_array[ 846 ] <= 16'hcb01;
mem_array[ 847 ] <= 16'hcb01;
mem_array[ 848 ] <= 16'hcb01;
mem_array[ 849 ] <= 16'hcb01;
mem_array[ 850 ] <= 16'hcb01;
mem_array[ 851 ] <= 16'hcb01;
mem_array[ 852 ] <= 16'hcb01;
mem_array[ 853 ] <= 16'hcb01;
mem_array[ 854 ] <= 16'hb241;
mem_array[ 855 ] <= 16'hb241;
mem_array[ 856 ] <= 16'hb241;
mem_array[ 857 ] <= 16'h9981;
mem_array[ 858 ] <= 16'h1;
mem_array[ 859 ] <= 16'h0;
mem_array[ 860 ] <= 16'h0;
mem_array[ 861 ] <= 16'h0;
mem_array[ 862 ] <= 16'h0;
mem_array[ 863 ] <= 16'h0;
mem_array[ 864 ] <= 16'h0;
mem_array[ 865 ] <= 16'h0;
mem_array[ 866 ] <= 16'h0;
mem_array[ 867 ] <= 16'h0;
mem_array[ 868 ] <= 16'h0;
mem_array[ 869 ] <= 16'h1;
mem_array[ 870 ] <= 16'h1;
mem_array[ 871 ] <= 16'h1;
mem_array[ 872 ] <= 16'h69c3;
mem_array[ 873 ] <= 16'hdbc5;
mem_array[ 874 ] <= 16'h1;
mem_array[ 875 ] <= 16'h9a41;
mem_array[ 876 ] <= 16'h5941;
mem_array[ 877 ] <= 16'h1;
mem_array[ 878 ] <= 16'h1;
mem_array[ 879 ] <= 16'h1;
mem_array[ 880 ] <= 16'h1;
mem_array[ 881 ] <= 16'hcb01;
mem_array[ 882 ] <= 16'hcb01;
mem_array[ 883 ] <= 16'hcb01;
mem_array[ 884 ] <= 16'hcb01;
mem_array[ 885 ] <= 16'hcb01;
mem_array[ 886 ] <= 16'hb241;
mem_array[ 887 ] <= 16'hb241;
mem_array[ 888 ] <= 16'h9981;
mem_array[ 889 ] <= 16'h1;
mem_array[ 890 ] <= 16'h0;
mem_array[ 891 ] <= 16'h0;
mem_array[ 892 ] <= 16'h0;
mem_array[ 893 ] <= 16'h0;
mem_array[ 894 ] <= 16'h0;
mem_array[ 895 ] <= 16'h0;
mem_array[ 896 ] <= 16'h0;
mem_array[ 897 ] <= 16'h0;
mem_array[ 898 ] <= 16'h0;
mem_array[ 899 ] <= 16'h0;
mem_array[ 900 ] <= 16'h0;
mem_array[ 901 ] <= 16'h0;
mem_array[ 902 ] <= 16'h1;
mem_array[ 903 ] <= 16'h1;
mem_array[ 904 ] <= 16'h1;
mem_array[ 905 ] <= 16'hcb01;
mem_array[ 906 ] <= 16'h1;
mem_array[ 907 ] <= 16'hcb01;
mem_array[ 908 ] <= 16'hcb01;
mem_array[ 909 ] <= 16'hcb01;
mem_array[ 910 ] <= 16'hcb01;
mem_array[ 911 ] <= 16'hcb01;
mem_array[ 912 ] <= 16'h1;
mem_array[ 913 ] <= 16'h1;
mem_array[ 914 ] <= 16'h1;
mem_array[ 915 ] <= 16'hcb01;
mem_array[ 916 ] <= 16'hb241;
mem_array[ 917 ] <= 16'hb241;
mem_array[ 918 ] <= 16'hb241;
mem_array[ 919 ] <= 16'h1;
mem_array[ 920 ] <= 16'h1;
mem_array[ 921 ] <= 16'h0;
mem_array[ 922 ] <= 16'h0;
mem_array[ 923 ] <= 16'h0;
mem_array[ 924 ] <= 16'h0;
mem_array[ 925 ] <= 16'h0;
mem_array[ 926 ] <= 16'h0;
mem_array[ 927 ] <= 16'h0;
mem_array[ 928 ] <= 16'h0;
mem_array[ 929 ] <= 16'h0;
mem_array[ 930 ] <= 16'h0;
mem_array[ 931 ] <= 16'h0;
mem_array[ 932 ] <= 16'h0;
mem_array[ 933 ] <= 16'h0;
mem_array[ 934 ] <= 16'h0;
mem_array[ 935 ] <= 16'h0;
mem_array[ 936 ] <= 16'h1;
mem_array[ 937 ] <= 16'h1;
mem_array[ 938 ] <= 16'h1;
mem_array[ 939 ] <= 16'h79c1;
mem_array[ 940 ] <= 16'hcb01;
mem_array[ 941 ] <= 16'hcb01;
mem_array[ 942 ] <= 16'hcb01;
mem_array[ 943 ] <= 16'hcb01;
mem_array[ 944 ] <= 16'hcb01;
mem_array[ 945 ] <= 16'hcb01;
mem_array[ 946 ] <= 16'hcb01;
mem_array[ 947 ] <= 16'h1;
mem_array[ 948 ] <= 16'h1;
mem_array[ 949 ] <= 16'h1;
mem_array[ 950 ] <= 16'h1;
mem_array[ 951 ] <= 16'h1;
mem_array[ 952 ] <= 16'h0;
mem_array[ 953 ] <= 16'h0;
mem_array[ 954 ] <= 16'h0;
mem_array[ 955 ] <= 16'h0;
mem_array[ 956 ] <= 16'h0;
mem_array[ 957 ] <= 16'h0;
mem_array[ 958 ] <= 16'h0;
mem_array[ 959 ] <= 16'h0;
mem_array[ 960 ] <= 16'h0;
mem_array[ 961 ] <= 16'h0;
mem_array[ 962 ] <= 16'h0;
mem_array[ 963 ] <= 16'h0;
mem_array[ 964 ] <= 16'h0;
mem_array[ 965 ] <= 16'h0;
mem_array[ 966 ] <= 16'h0;
mem_array[ 967 ] <= 16'h0;
mem_array[ 968 ] <= 16'h0;
mem_array[ 969 ] <= 16'h0;
mem_array[ 970 ] <= 16'h1;
mem_array[ 971 ] <= 16'h1;
mem_array[ 972 ] <= 16'h1;
mem_array[ 973 ] <= 16'h1;
mem_array[ 974 ] <= 16'h1;
mem_array[ 975 ] <= 16'h1;
mem_array[ 976 ] <= 16'h1;
mem_array[ 977 ] <= 16'h1;
mem_array[ 978 ] <= 16'h1;
mem_array[ 979 ] <= 16'h1;
mem_array[ 980 ] <= 16'h1;
mem_array[ 981 ] <= 16'h1;
mem_array[ 982 ] <= 16'h0;
mem_array[ 983 ] <= 16'h0;
mem_array[ 984 ] <= 16'h0;
mem_array[ 985 ] <= 16'h0;
mem_array[ 986 ] <= 16'h0;
mem_array[ 987 ] <= 16'h0;
mem_array[ 988 ] <= 16'h0;
mem_array[ 989 ] <= 16'h0;
mem_array[ 990 ] <= 16'h0;
mem_array[ 991 ] <= 16'h0;
mem_array[ 992 ] <= 16'h0;
mem_array[ 993 ] <= 16'h0;
mem_array[ 994 ] <= 16'h0;
mem_array[ 995 ] <= 16'h0;
mem_array[ 996 ] <= 16'h0;
mem_array[ 997 ] <= 16'h0;
mem_array[ 998 ] <= 16'h0;
mem_array[ 999 ] <= 16'h0;
mem_array[ 1000 ] <= 16'h0;
mem_array[ 1001 ] <= 16'h0;
mem_array[ 1002 ] <= 16'h0;
mem_array[ 1003 ] <= 16'h0;
mem_array[ 1004 ] <= 16'h0;
mem_array[ 1005 ] <= 16'h0;
mem_array[ 1006 ] <= 16'h1;
mem_array[ 1007 ] <= 16'h1;
mem_array[ 1008 ] <= 16'h1;
mem_array[ 1009 ] <= 16'h1;
mem_array[ 1010 ] <= 16'h7bdf;
mem_array[ 1011 ] <= 16'h0;
mem_array[ 1012 ] <= 16'h0;
mem_array[ 1013 ] <= 16'h0;
mem_array[ 1014 ] <= 16'h0;
mem_array[ 1015 ] <= 16'h0;
mem_array[ 1016 ] <= 16'h0;
mem_array[ 1017 ] <= 16'h0;
mem_array[ 1018 ] <= 16'h0;
mem_array[ 1019 ] <= 16'h0;
mem_array[ 1020 ] <= 16'h0;
mem_array[ 1021 ] <= 16'h0;
mem_array[ 1022 ] <= 16'h0;
mem_array[ 1023 ] <= 16'h0;


			
			for (integer i = 1024; i <= size - 1; i = i + 1)		// Assign the rest of the memory to 0
			begin
				mem_array[i] <= 16'h0;
			end
		end
		else if (~CE && ~WE)
		begin
            if(~UB)
			    mem_array[A[10:0]][15:8] <= I_O[15:8];   // A(15 downto X+1): X must
														// be the same as above
		    if(~LB)
			    mem_array[A[10:0]][7:0] <= I_O[7:0];     // A(X downto 0): X
		end                                             // must be the same as above

   end
	  
   assign I_O = I_O_wire;
	  
endmodule