/**
 * SpriteDrawer.sv
 * 
 * A state machine that read sprite data from sram given the current vga coordinate
 * 
 */


module SpirteDrawer(
	input logic[19:0] A,
	input logic[9:0] DrawX, DrawY,
	
	output logic[7:0] R, G, B 
)



endmodule 